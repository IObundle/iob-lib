   //General interface signals (do not remove indentation)
   //START_IO_TABLE gen
   `IOB_INPUT(clk,          1), //System clock input
   `IOB_INPUT(rst,          1)  //System reset, asynchronous and active high
