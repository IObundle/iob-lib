   //General interface signals (do not remove indentation)
   //START_IO_TABLE gen
   `INPUT(clk,          1), //System clock input
   `INPUT(rst,          1)  //System reset, asynchronous and active high
