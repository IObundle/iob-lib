   //General Interface Signals (do not remove indentation)
   //START_IO_TABLE gen
   input [1-1:0] clk_i, //V2TEX_IO System clock.
   input [1-1:0] cke_i,  //V2TEX_IO System clock enable.
   input [1-1:0] arst_i  //V2TEX_IO System reset, asynchronous and active high.
