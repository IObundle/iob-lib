`define BAUD 115200
`define FREQ 100000000
`define DDR_DATA_W 32
`define DDR_ADDR_W 30
`define MEM_ADDR_W 24
`define XILINX 1
