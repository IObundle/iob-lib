      .clk_i(clk_i),
      .arst_i(arst_i)
