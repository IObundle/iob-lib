`timescale 1ns/1ps

`include "iob_lib.vh"

module iob_fifo_async
  #(parameter
    W_DATA_W = 0,
    R_DATA_W = 0,
    ADDR_W = 0, //higher ADDR_W lower DATA_W
    //determine W_ADDR_W and R_ADDR_W
   MAXDATA_W = `IOB_MAX(W_DATA_W, R_DATA_W),
   MINDATA_W = `IOB_MIN(W_DATA_W, R_DATA_W),
   R = MAXDATA_W/MINDATA_W,
   ADDR_W_DIFF = $clog2(R),
   MINADDR_W = ADDR_W-$clog2(R),//lower ADDR_W (higher DATA_W)
   W_ADDR_W = (W_DATA_W == MAXDATA_W) ? MINADDR_W : ADDR_W,
   R_ADDR_W = (R_DATA_W == MAXDATA_W) ? MINADDR_W : ADDR_W
    )
   (
      
   //memory write port
   `IOB_OUTPUT(ext_mem_w_clk_o, 1),
   `IOB_OUTPUT(ext_mem_w_en_o, 1),
   `IOB_OUTPUT(ext_mem_w_addr_o, W_ADDR_W),
   `IOB_OUTPUT(ext_mem_w_data_o, W_DATA_W),
   //memory read port
   `IOB_OUTPUT(ext_mem_r_clk_o, 1),
   `IOB_OUTPUT(ext_mem_r_en_o, 1),
   `IOB_OUTPUT(ext_mem_r_addr_o, R_ADDR_W),
   `IOB_INPUT(ext_mem_r_data_i, R_DATA_W),
    
    //read port
    input                 r_clk_i,
    input                 r_arst_i,
    input                 r_cke_i,
    input                 r_rst_i,
    input                 r_en_i,
    output [R_DATA_W-1:0] r_data_o,
    output                r_empty_o,
    output                r_full_o,
    output [ADDR_W:0]     r_level_o,

    //write port
    input                 w_clk_i,
    input                 w_arst_i,
    input                 w_cke_i,
    input                 w_rst_i,
    input                 w_en_i,
    input [W_DATA_W-1:0]  w_data_i,
    output                w_empty_o,
    output                w_full_o,
    output [ADDR_W:0]     w_level_o

    );

   localparam [ADDR_W:0] FIFO_SIZE = (1'b1 << ADDR_W); //in bytes

   //binary read addresses on both domains
   wire [R_ADDR_W:0]        r_raddr_bin;
   wire [R_ADDR_W:0]        w_raddr_bin;
   wire [W_ADDR_W:0]        r_waddr_bin;
   wire [W_ADDR_W:0]        w_waddr_bin;

   //normalized binary addresses (for narrower data side)
   wire [ADDR_W:0]          r_raddr_bin_n;
   wire [ADDR_W:0]          r_waddr_bin_n;
   wire [ADDR_W:0]          w_waddr_bin_n;
   wire [ADDR_W:0]          w_raddr_bin_n;

   //assign according to assymetry type
   localparam [ADDR_W-1:0] w_incr = (W_DATA_W > R_DATA_W) ? 1'b1 << ADDR_W_DIFF : 1'b1 ;
   localparam [ADDR_W-1:0] r_incr = (R_DATA_W > W_DATA_W) ? 1'b1 << ADDR_W_DIFF : 1'b1 ;
   
   generate
      if (W_DATA_W > R_DATA_W) begin
         assign w_waddr_bin_n = w_waddr_bin<<ADDR_W_DIFF;
         assign w_raddr_bin_n = w_raddr_bin;
         assign r_raddr_bin_n = r_raddr_bin;
         assign r_waddr_bin_n = r_waddr_bin<<ADDR_W_DIFF;
      end else if (R_DATA_W > W_DATA_W) begin
         assign w_waddr_bin_n = w_waddr_bin;
         assign w_raddr_bin_n = w_raddr_bin<<ADDR_W_DIFF;
         assign r_raddr_bin_n = r_raddr_bin<<ADDR_W_DIFF;
         assign r_waddr_bin_n = r_waddr_bin;
      end else begin
         assign w_raddr_bin_n = w_raddr_bin;
         assign w_waddr_bin_n = w_waddr_bin;
         assign r_waddr_bin_n = r_waddr_bin;
         assign r_raddr_bin_n = r_raddr_bin;
      end
   endgenerate


   //sync write gray address to read domain
   wire [W_ADDR_W:0]        w_waddr_gray;
   wire [W_ADDR_W:0]        r_waddr_gray;
   iob_sync
     #(
       .DATA_W(W_ADDR_W+1),
       .RST_VAL(0)
       )
   w_waddr_gray_sync0
     (
      .clk_i    (r_clk_i),
      .arst_i   (r_arst_i),
      .cke_i    (r_cke_i),
      .signal_i (w_waddr_gray),
      .signal_o (r_waddr_gray)
      );

   //sync read gray address to write domain
   wire [R_ADDR_W:0]        r_raddr_gray;
   wire [R_ADDR_W:0]        w_raddr_gray;
   iob_sync
     #(
       .DATA_W(R_ADDR_W+1),
       .RST_VAL(0)
       )
   r_raddr_gray_sync0
     (
      .clk_i    (w_clk_i),
      .arst_i   (w_arst_i),
      .cke_i    (w_cke_i),
      .signal_i (r_raddr_gray),
      .signal_o (w_raddr_gray)
      );


   //READ DOMAIN FIFO LEVEL
   `IOB_WIRE(r_level_int, (ADDR_W+2))
   assign r_level_int = r_waddr_bin_n - r_raddr_bin_n;
   assign r_level_o = r_level_int[0+:(ADDR_W+1)];
   
   //READ DOMAIN EMPTY AND FULL FLAGS
   assign r_empty_o = (r_level_int < {2'd0, r_incr});
   `IOB_WIRE(r_full_limit, (ADDR_W+2))
   assign r_full_limit = FIFO_SIZE-{2'd0, r_incr};
   assign r_full_o = (r_level_int > r_full_limit);

   //WRITE DOMAIN FIFO LEVEL
   `IOB_WIRE(w_level_int, (ADDR_W+2))
   assign w_level_int = w_waddr_bin_n - w_raddr_bin_n;
   assign w_level_o = w_level_int[0+:(ADDR_W+1)];
 
   //WRITE DOMAIN EMPTY AND FULL FLAGS
   assign w_empty_o = (w_level_int < {2'd0, w_incr});
   `IOB_WIRE(w_full_limit, (ADDR_W+2))
   assign w_full_limit = FIFO_SIZE-{2'd0, w_incr};
   assign w_full_o = (w_level_int > w_full_limit);

   
   //read address gray code counter
   wire r_en_int  = (r_en_i & (~r_empty_o));
   iob_gray_counter
     #(
       .W(R_ADDR_W+1)
       )
   r_raddr_gray_counter
     (
      .clk_i  (r_clk_i),
      .arst_i (r_arst_i),
      .cke_i  (r_cke_i),
      .rst_i  (r_rst_i),
      .en_i   (r_en_int),
      .data_o (r_raddr_gray)
      );

   //write address gray code counter
   wire w_en_int = (w_en_i & (~w_full_o));
   iob_gray_counter
     #(
       .W(W_ADDR_W+1)
       )
   w_waddr_gray_counter
     (
      .clk_i  (w_clk_i),
      .arst_i (w_arst_i),
      .cke_i  (w_cke_i),
      .rst_i  (w_rst_i),
      .en_i   (w_en_int),
      .data_o (w_waddr_gray)
      );

   //convert gray read address to binary
   iob_gray2bin
     #(
       .DATA_W(R_ADDR_W+1)
       )
   gray2bin_r_raddr
     (
      .gr_i  (r_raddr_gray),
      .bin_o (r_raddr_bin)
      );

   //convert synced gray write address to binary
   iob_gray2bin
     #(
       .DATA_W(W_ADDR_W+1)
       )
   gray2bin_r_raddr_sync
     (
      .gr_i  (r_waddr_gray),
      .bin_o (r_waddr_bin)
      );

   //convert gray write address to binary
   iob_gray2bin
     #(
       .DATA_W(W_ADDR_W+1)
       )
   gray2bin_w_waddr
     (
      .gr_i  (w_waddr_gray),
      .bin_o (w_waddr_bin)
      );

   //convert synced gray read address to binary
   iob_gray2bin
     #(
       .DATA_W(R_ADDR_W+1)
       )
   gray2bin_w_raddr_sync
     (
      .gr_i  (w_raddr_gray),
      .bin_o (w_raddr_bin)
      );

   // FIFO memory
   assign ext_mem_w_clk_o = w_clk_i;
   assign ext_mem_w_en_o = w_en_int;
   assign ext_mem_w_addr_o = w_waddr_bin[W_ADDR_W-1:0];
   assign ext_mem_w_data_o = w_data_i;
   assign ext_mem_r_clk_o = r_clk_i;
   assign ext_mem_r_en_o = r_en_int;
   assign ext_mem_r_addr_o = r_raddr_bin[R_ADDR_W-1:0];
   assign r_data_o = ext_mem_r_data_i;

endmodule
