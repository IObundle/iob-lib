//General interface signals (do not remove indentation)
    //START_TABLE gen_if
   `INPUT(clk,          1), //System clock input
   `INPUT(rst,          1) //System reset, asynchronous and active high
