.iob_avalid_o(iob_avalid), //Request valid.
.iob_addr_o(iob_addr), //Address.
.iob_wdata_o(iob_wdata), //Write data.
.iob_wstrb_o(iob_wstrb), //Write strobe.
.iob_rvalid_nxt_i(iob_rvalid_nxt), //Read data valid.
.iob_rdata_i(iob_rdata), //Read data.
.iob_ready_nxt_i(iob_ready_nxt), //Interface ready.
