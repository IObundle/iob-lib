      .valid(valid),
      .ready(ready),
      .addr(addr),
      .wdata(wdata),
      .wstrb(wstrb),
      .rvalid(rvalid),
      .rdata(rdata),
