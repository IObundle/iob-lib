      .clk_i(clk_i),
      .en_i(en_i),
      .arst_i(arst_i)
