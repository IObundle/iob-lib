      .clk_i(clk_i),
      .rst_i(rst_i)
