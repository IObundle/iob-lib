      .clk_i(clk_i),
      .cke_i(cke_i),
      .arst_i(arst_i)
