`timescale 1ns / 1ps

`include "iob_lib.vh"

module axil2iob
  #(
    parameter AXIL_ADDR_W = 32,     // AXI Lite address bus width in bits
    parameter AXIL_DATA_W = 32,     // AXI Lite data bus width in bits
    parameter ADDR_W = AXIL_ADDR_W, // IOb address bus width in bits
    parameter DATA_W = AXIL_DATA_W  // IOb data bus width in bits
    )
   (
    // AXI4 Lite slave interface
`include "axil_s_port.vh"

    // IOb master interface
`include "iob_m_port.vh"

    // Global signals
`include "iob_clkrst_port.vh"
    );

   //
   // COMPUTE AXIL OUTPUTS
   //
   
   // write address
   assign axil_awready_o = iob_ready_i;

   // write
   assign axil_wready_o = iob_ready_i;

   // write response
   assign axil_bresp_o = 2'b0;
   assign axil_bvalid_o = 1'b1;

   // read address
   assign axil_arready_o = iob_ready_i;

   // read
   assign axil_rdata_o = iob_rdata_i;
   assign axil_rresp_o = 2'b0;
   assign axil_rvalid_o = iob_rvalid_i;

   //
   // COMPUTE IOb OUTPUTS
   //
   assign iob_valid_o = axil_awvalid_i | axil_wvalid_i | axil_arvalid_i;
   assign iob_addr_o  = axil_awvalid_i? axil_awaddr_i: axil_araddr_i;
   assign iob_wdata_o = axil_wdata_i;
   assign iob_wstrb_o = axil_wvalid_i? axil_wstrb_i: {DATA_W/8{1'b0}};

endmodule
