      .valid_o  (valid_i),
      .ready_i  (ready_o),
      .addr_o   (addr_i),
      .wdata_o  (wdata_i),
      .wstrb_o  (wstrb_i),
      .rvalid_i (rvalid_o),
      .rdata_i  (rdata_o),
