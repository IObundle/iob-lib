   //General Interface Signals (do not remove indentation)
   //START_IO_TABLE gen
   `IOB_INPUT(clk_i,          1), //V2TEX_IO System clock.
   `IOB_INPUT(cke_i,          1),  //V2TEX_IO System clock enable.
   `IOB_INPUT(arst_i,         1)  //V2TEX_IO System reset, asynchronous and active high.
