      .valid_i  (valid_o),
      .ready_o  (ready_i),
      .addr_i   (addr_o),
      .wdata_i  (wdata_o),
      .wstrb_i  (wstrb_o),
      .rvalid_o (rvalid_i),
      .rdata_o  (rdata_i),
